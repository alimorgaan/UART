module baud_test ();


baud


endmodule